module if_id(
    input clk,
    input rst_n,
    // from instruction fetch

    // to instruction decode

);


endmodule